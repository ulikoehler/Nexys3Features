../../util/clkdiv_rst/src/clkdiv_rst.vhd